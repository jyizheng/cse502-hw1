
`ifndef _GPR_SVH_
`define _GPR_SVH_ 1


/* RFLAGS fields */

`define RF_IMPL_MSB	31
`define RF_IMPL_LSB	28
`define RF_VER_MSB	27
`define RF_VER_LSB	24
`define RF_ICC_MSB	23
`define RF_ICC_LSB	20
`define RF_N	23
`define RF_Z	22
`define RF_V	21
`define RF_C	20
`define RF_RESV_MSB	19
`define RF_RESV_LSB	14
`define RF_EC	13
`define RF_EF	12
`define RF_PIL_MSB	11
`define RF_PIL_LSB	8
`define RF_S	7
`define RF_PS	6
`define RF_ET	5
`define RF_CWP_MSB	4
`define RF_CWP_LSB	0


`endif

/* vim: set ts=4 sw=0 tw=0 noet : */
