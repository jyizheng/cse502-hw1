`ifndef _GLOBAL_SVH_
`define _GLOBAL_SVH_ 1

`define REG_TOTAL_NUM	32

`define REG_WIN_NUM	144
`define REG_GLB_NUM	8
`define REG_IN_NUM	8
`define REG_LOCAL_NUM	8
`define REG_OUT_NUM	8


`endif

